* NGSPICE file created from dec_to_bin.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

.subckt dec_to_bin vdd gnd decimal[0] decimal[1] decimal[2] decimal[3] decimal[4]
+ decimal[5] decimal[6] decimal[7] octal[0] octal[1] octal[2] octal[3] octal[4] octal[5]
+ octal[6] octal[7]
XFILL_0_0_0 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XFILL_0_0_2 gnd vdd FILL
XBUFX2_1 decimal[0] gnd octal[0] vdd BUFX2
XBUFX2_2 decimal[1] gnd octal[1] vdd BUFX2
XBUFX2_3 decimal[2] gnd octal[2] vdd BUFX2
XBUFX2_4 decimal[3] gnd octal[3] vdd BUFX2
XBUFX2_5 decimal[4] gnd octal[4] vdd BUFX2
XFILL_0_1_0 gnd vdd FILL
XBUFX2_6 decimal[5] gnd octal[5] vdd BUFX2
XFILL_0_1_1 gnd vdd FILL
XBUFX2_7 decimal[6] gnd octal[6] vdd BUFX2
XFILL_0_1_2 gnd vdd FILL
XBUFX2_8 decimal[7] gnd octal[7] vdd BUFX2
.ends

