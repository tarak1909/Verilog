VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dec_to_hex
  CLASS BLOCK ;
  FOREIGN dec_to_hex ;
  ORIGIN 1.900 0.000 ;
  SIZE 53.400 BY 26.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 2.800 1.600 3.600 9.000 ;
        RECT 7.600 1.600 8.400 9.000 ;
        RECT 17.200 1.600 18.000 9.000 ;
        RECT 22.000 1.600 22.800 9.000 ;
        RECT 26.800 1.600 27.600 9.000 ;
        RECT 31.600 1.600 32.400 9.000 ;
        RECT 41.200 1.600 42.000 9.000 ;
        RECT 46.000 1.600 46.800 9.000 ;
        RECT 0.400 0.400 49.200 1.600 ;
      LAYER via1 ;
        RECT 11.000 0.600 11.800 1.400 ;
        RECT 12.400 0.600 13.200 1.400 ;
        RECT 13.800 0.600 14.600 1.400 ;
      LAYER metal2 ;
        RECT 10.400 0.600 15.200 1.400 ;
      LAYER via2 ;
        RECT 11.000 0.600 11.800 1.400 ;
        RECT 12.400 0.600 13.200 1.400 ;
        RECT 13.800 0.600 14.600 1.400 ;
      LAYER metal3 ;
        RECT 10.400 0.400 15.200 1.600 ;
      LAYER via3 ;
        RECT 10.800 0.600 11.600 1.400 ;
        RECT 12.400 0.600 13.200 1.400 ;
        RECT 14.000 0.600 14.800 1.400 ;
      LAYER metal4 ;
        RECT 10.400 0.000 15.200 24.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.400 20.400 49.200 21.600 ;
        RECT 2.800 15.800 3.600 20.400 ;
        RECT 7.600 15.800 8.400 20.400 ;
        RECT 17.200 15.800 18.000 20.400 ;
        RECT 22.000 15.800 22.800 20.400 ;
        RECT 26.800 15.800 27.600 20.400 ;
        RECT 31.600 15.800 32.400 20.400 ;
        RECT 41.200 15.800 42.000 20.400 ;
        RECT 46.000 15.800 46.800 20.400 ;
      LAYER via1 ;
        RECT 35.000 20.600 35.800 21.400 ;
        RECT 36.400 20.600 37.200 21.400 ;
        RECT 37.800 20.600 38.600 21.400 ;
      LAYER metal2 ;
        RECT 34.400 20.600 39.200 21.400 ;
      LAYER via2 ;
        RECT 35.000 20.600 35.800 21.400 ;
        RECT 36.400 20.600 37.200 21.400 ;
        RECT 37.800 20.600 38.600 21.400 ;
      LAYER metal3 ;
        RECT 34.400 20.400 39.200 21.600 ;
      LAYER via3 ;
        RECT 34.800 20.600 35.600 21.400 ;
        RECT 36.400 20.600 37.200 21.400 ;
        RECT 38.000 20.600 38.800 21.400 ;
      LAYER metal4 ;
        RECT 34.400 0.000 39.200 24.000 ;
    END
  END gnd
  PIN decimal[0]
    PORT
      LAYER metal1 ;
        RECT 10.800 12.300 11.600 12.400 ;
        RECT 15.600 12.300 16.400 13.200 ;
        RECT 10.800 11.700 16.400 12.300 ;
        RECT 10.800 11.600 11.600 11.700 ;
        RECT 15.600 11.600 16.400 11.700 ;
      LAYER metal2 ;
        RECT 7.700 20.400 8.300 24.300 ;
        RECT 7.600 19.600 8.400 20.400 ;
        RECT 10.800 19.600 11.600 20.400 ;
        RECT 10.900 12.400 11.500 19.600 ;
        RECT 10.800 11.600 11.600 12.400 ;
      LAYER metal3 ;
        RECT 7.600 20.300 8.400 20.400 ;
        RECT 10.800 20.300 11.600 20.400 ;
        RECT 7.600 19.700 11.600 20.300 ;
        RECT 7.600 19.600 8.400 19.700 ;
        RECT 10.800 19.600 11.600 19.700 ;
    END
  END decimal[0]
  PIN decimal[1]
    PORT
      LAYER metal1 ;
        RECT 39.600 11.600 40.400 13.200 ;
      LAYER metal2 ;
        RECT 39.700 25.700 43.500 26.300 ;
        RECT 39.700 24.300 40.300 25.700 ;
        RECT 36.500 23.700 40.300 24.300 ;
        RECT 42.900 20.400 43.500 25.700 ;
        RECT 42.800 19.600 43.600 20.400 ;
        RECT 39.600 11.600 40.400 12.400 ;
        RECT 39.700 10.400 40.300 11.600 ;
        RECT 39.600 9.600 40.400 10.400 ;
      LAYER metal3 ;
        RECT 42.800 19.600 43.600 20.400 ;
        RECT 39.600 10.300 40.400 10.400 ;
        RECT 42.800 10.300 43.600 10.400 ;
        RECT 39.600 9.700 43.600 10.300 ;
        RECT 39.600 9.600 40.400 9.700 ;
        RECT 42.800 9.600 43.600 9.700 ;
      LAYER metal4 ;
        RECT 42.600 9.400 43.800 20.600 ;
    END
  END decimal[1]
  PIN decimal[2]
    PORT
      LAYER metal1 ;
        RECT 23.600 11.600 24.400 13.200 ;
      LAYER metal2 ;
        RECT 23.700 23.700 25.900 24.300 ;
        RECT 23.700 12.400 24.300 23.700 ;
        RECT 23.600 11.600 24.400 12.400 ;
    END
  END decimal[2]
  PIN decimal[3]
    PORT
      LAYER metal1 ;
        RECT 44.400 11.600 45.200 13.200 ;
      LAYER metal2 ;
        RECT 41.300 14.400 41.900 24.300 ;
        RECT 41.200 13.600 42.000 14.400 ;
        RECT 44.400 13.600 45.200 14.400 ;
        RECT 44.500 12.400 45.100 13.600 ;
        RECT 44.400 11.600 45.200 12.400 ;
      LAYER metal3 ;
        RECT 41.200 14.300 42.000 14.400 ;
        RECT 44.400 14.300 45.200 14.400 ;
        RECT 41.200 13.700 45.200 14.300 ;
        RECT 41.200 13.600 42.000 13.700 ;
        RECT 44.400 13.600 45.200 13.700 ;
    END
  END decimal[3]
  PIN decimal[4]
    PORT
      LAYER metal1 ;
        RECT 4.400 11.600 5.200 13.200 ;
      LAYER metal2 ;
        RECT 2.800 19.600 3.600 20.400 ;
        RECT 2.900 16.300 3.500 19.600 ;
        RECT 2.900 15.700 5.100 16.300 ;
        RECT 4.500 12.400 5.100 15.700 ;
        RECT 4.400 11.600 5.200 12.400 ;
      LAYER metal3 ;
        RECT 2.800 20.300 3.600 20.400 ;
        RECT -1.900 19.700 3.600 20.300 ;
        RECT 2.800 19.600 3.600 19.700 ;
    END
  END decimal[4]
  PIN decimal[5]
    PORT
      LAYER metal1 ;
        RECT 25.200 11.600 26.000 13.200 ;
      LAYER metal2 ;
        RECT 28.500 20.400 29.100 24.300 ;
        RECT 25.200 19.600 26.000 20.400 ;
        RECT 28.400 19.600 29.200 20.400 ;
        RECT 25.300 12.400 25.900 19.600 ;
        RECT 25.200 11.600 26.000 12.400 ;
      LAYER metal3 ;
        RECT 25.200 20.300 26.000 20.400 ;
        RECT 28.400 20.300 29.200 20.400 ;
        RECT 25.200 19.700 29.200 20.300 ;
        RECT 25.200 19.600 26.000 19.700 ;
        RECT 28.400 19.600 29.200 19.700 ;
    END
  END decimal[5]
  PIN decimal[6]
    PORT
      LAYER metal1 ;
        RECT 9.200 11.600 10.000 13.200 ;
      LAYER metal2 ;
        RECT 4.500 18.400 5.100 24.300 ;
        RECT 4.400 17.600 5.200 18.400 ;
        RECT 9.200 17.600 10.000 18.400 ;
        RECT 9.300 12.400 9.900 17.600 ;
        RECT 9.200 11.600 10.000 12.400 ;
      LAYER metal3 ;
        RECT 4.400 18.300 5.200 18.400 ;
        RECT 9.200 18.300 10.000 18.400 ;
        RECT 4.400 17.700 10.000 18.300 ;
        RECT 4.400 17.600 5.200 17.700 ;
        RECT 9.200 17.600 10.000 17.700 ;
    END
  END decimal[6]
  PIN decimal[7]
    PORT
      LAYER metal1 ;
        RECT 30.000 11.600 30.800 13.200 ;
      LAYER metal2 ;
        RECT 46.000 19.600 46.800 20.400 ;
        RECT 46.100 16.400 46.700 19.600 ;
        RECT 30.000 15.600 30.800 16.400 ;
        RECT 46.000 15.600 46.800 16.400 ;
        RECT 30.100 12.400 30.700 15.600 ;
        RECT 30.000 11.600 30.800 12.400 ;
      LAYER metal3 ;
        RECT 46.000 20.300 46.800 20.400 ;
        RECT 46.000 19.700 51.500 20.300 ;
        RECT 46.000 19.600 46.800 19.700 ;
        RECT 30.000 16.300 30.800 16.400 ;
        RECT 46.000 16.300 46.800 16.400 ;
        RECT 30.000 15.700 46.800 16.300 ;
        RECT 30.000 15.600 30.800 15.700 ;
        RECT 46.000 15.600 46.800 15.700 ;
    END
  END decimal[7]
  PIN hex[0]
    PORT
      LAYER metal1 ;
        RECT 18.800 12.400 19.600 19.800 ;
        RECT 19.000 10.200 19.600 12.400 ;
        RECT 18.800 2.200 19.600 10.200 ;
      LAYER via1 ;
        RECT 18.800 17.600 19.600 18.400 ;
      LAYER metal2 ;
        RECT 12.500 20.400 13.100 24.300 ;
        RECT 12.400 19.600 13.200 20.400 ;
        RECT 18.800 19.600 19.600 20.400 ;
        RECT 18.900 18.400 19.500 19.600 ;
        RECT 18.800 17.600 19.600 18.400 ;
      LAYER metal3 ;
        RECT 12.400 20.300 13.200 20.400 ;
        RECT 18.800 20.300 19.600 20.400 ;
        RECT 12.400 19.700 19.600 20.300 ;
        RECT 12.400 19.600 13.200 19.700 ;
        RECT 18.800 19.600 19.600 19.700 ;
    END
  END hex[0]
  PIN hex[1]
    PORT
      LAYER metal1 ;
        RECT 42.800 12.400 43.600 19.800 ;
        RECT 43.000 10.200 43.600 12.400 ;
        RECT 42.800 2.200 43.600 10.200 ;
      LAYER via1 ;
        RECT 42.800 13.600 43.600 14.400 ;
      LAYER metal2 ;
        RECT 42.800 13.600 43.600 14.400 ;
        RECT 42.900 12.400 43.500 13.600 ;
        RECT 42.800 11.600 43.600 12.400 ;
      LAYER metal3 ;
        RECT 42.800 12.300 43.600 12.400 ;
        RECT 42.800 11.700 51.500 12.300 ;
        RECT 42.800 11.600 43.600 11.700 ;
    END
  END hex[1]
  PIN hex[2]
    PORT
      LAYER metal1 ;
        RECT 20.400 12.400 21.200 19.800 ;
        RECT 20.400 10.200 21.000 12.400 ;
        RECT 20.400 2.200 21.200 10.200 ;
      LAYER via1 ;
        RECT 20.400 17.600 21.200 18.400 ;
      LAYER metal2 ;
        RECT 15.700 18.400 16.300 24.300 ;
        RECT 15.600 17.600 16.400 18.400 ;
        RECT 20.400 17.600 21.200 18.400 ;
      LAYER metal3 ;
        RECT 15.600 18.300 16.400 18.400 ;
        RECT 20.400 18.300 21.200 18.400 ;
        RECT 15.600 17.700 21.200 18.300 ;
        RECT 15.600 17.600 16.400 17.700 ;
        RECT 20.400 17.600 21.200 17.700 ;
    END
  END hex[2]
  PIN hex[3]
    PORT
      LAYER metal1 ;
        RECT 47.600 12.400 48.400 19.800 ;
        RECT 47.800 10.200 48.400 12.400 ;
        RECT 47.600 2.200 48.400 10.200 ;
      LAYER via1 ;
        RECT 47.600 17.600 48.400 18.400 ;
      LAYER metal2 ;
        RECT 47.700 23.700 49.900 24.300 ;
        RECT 47.700 18.400 48.300 23.700 ;
        RECT 47.600 17.600 48.400 18.400 ;
    END
  END hex[3]
  PIN hex[4]
    PORT
      LAYER metal1 ;
        RECT 1.200 12.400 2.000 19.800 ;
        RECT 1.200 10.200 1.800 12.400 ;
        RECT 1.200 2.200 2.000 10.200 ;
      LAYER via1 ;
        RECT 1.200 15.600 2.000 16.400 ;
      LAYER metal2 ;
        RECT 1.200 15.600 2.000 16.400 ;
      LAYER metal3 ;
        RECT 1.200 16.300 2.000 16.400 ;
        RECT -1.900 15.700 2.000 16.300 ;
        RECT 1.200 15.600 2.000 15.700 ;
    END
  END hex[4]
  PIN hex[5]
    PORT
      LAYER metal1 ;
        RECT 28.400 12.400 29.200 19.800 ;
        RECT 28.600 10.200 29.200 12.400 ;
        RECT 28.400 2.200 29.200 10.200 ;
      LAYER via1 ;
        RECT 28.400 17.600 29.200 18.400 ;
      LAYER metal2 ;
        RECT 31.700 23.700 33.900 24.300 ;
        RECT 31.700 18.400 32.300 23.700 ;
        RECT 28.400 17.600 29.200 18.400 ;
        RECT 31.600 17.600 32.400 18.400 ;
      LAYER metal3 ;
        RECT 28.400 18.300 29.200 18.400 ;
        RECT 31.600 18.300 32.400 18.400 ;
        RECT 28.400 17.700 32.400 18.300 ;
        RECT 28.400 17.600 29.200 17.700 ;
        RECT 31.600 17.600 32.400 17.700 ;
    END
  END hex[5]
  PIN hex[6]
    PORT
      LAYER metal1 ;
        RECT 6.000 12.400 6.800 19.800 ;
        RECT 6.000 10.200 6.600 12.400 ;
        RECT 6.000 2.200 6.800 10.200 ;
      LAYER via1 ;
        RECT 6.000 13.600 6.800 14.400 ;
      LAYER metal2 ;
        RECT 6.000 13.600 6.800 14.400 ;
        RECT 6.100 12.400 6.700 13.600 ;
        RECT 6.000 11.600 6.800 12.400 ;
      LAYER metal3 ;
        RECT 6.000 12.300 6.800 12.400 ;
        RECT -1.900 11.700 6.800 12.300 ;
        RECT 6.000 11.600 6.800 11.700 ;
    END
  END hex[6]
  PIN hex[7]
    PORT
      LAYER metal1 ;
        RECT 33.200 18.300 34.000 19.800 ;
        RECT 38.000 18.300 38.800 18.400 ;
        RECT 33.200 17.700 38.800 18.300 ;
        RECT 33.200 12.400 34.000 17.700 ;
        RECT 38.000 17.600 38.800 17.700 ;
        RECT 33.400 10.200 34.000 12.400 ;
        RECT 33.200 2.200 34.000 10.200 ;
      LAYER metal2 ;
        RECT 38.000 17.600 38.800 18.400 ;
      LAYER metal3 ;
        RECT 38.000 18.300 38.800 18.400 ;
        RECT 38.000 17.700 51.500 18.300 ;
        RECT 38.000 17.600 38.800 17.700 ;
        RECT 50.900 15.700 51.500 17.700 ;
    END
  END hex[7]
  OBS
      LAYER metal1 ;
        RECT 4.400 15.200 5.200 19.800 ;
        RECT 9.200 15.200 10.000 19.800 ;
        RECT 3.000 14.600 5.200 15.200 ;
        RECT 7.800 14.600 10.000 15.200 ;
        RECT 15.600 15.200 16.400 19.800 ;
        RECT 23.600 15.200 24.400 19.800 ;
        RECT 15.600 14.600 17.800 15.200 ;
        RECT 3.000 11.600 3.600 14.600 ;
        RECT 7.800 11.600 8.400 14.600 ;
        RECT 2.400 10.800 3.600 11.600 ;
        RECT 7.200 10.800 8.400 11.600 ;
        RECT 3.000 10.200 3.600 10.800 ;
        RECT 7.800 10.200 8.400 10.800 ;
        RECT 17.200 11.600 17.800 14.600 ;
        RECT 22.200 14.600 24.400 15.200 ;
        RECT 25.200 15.200 26.000 19.800 ;
        RECT 30.000 15.200 30.800 19.800 ;
        RECT 39.600 15.200 40.400 19.800 ;
        RECT 44.400 15.200 45.200 19.800 ;
        RECT 25.200 14.600 27.400 15.200 ;
        RECT 30.000 14.600 32.200 15.200 ;
        RECT 39.600 14.600 41.800 15.200 ;
        RECT 44.400 14.600 46.600 15.200 ;
        RECT 22.200 11.600 22.800 14.600 ;
        RECT 17.200 10.800 18.400 11.600 ;
        RECT 21.600 10.800 22.800 11.600 ;
        RECT 17.200 10.200 17.800 10.800 ;
        RECT 3.000 9.600 5.200 10.200 ;
        RECT 7.800 9.600 10.000 10.200 ;
        RECT 4.400 2.200 5.200 9.600 ;
        RECT 9.200 2.200 10.000 9.600 ;
        RECT 15.600 9.600 17.800 10.200 ;
        RECT 22.200 10.200 22.800 10.800 ;
        RECT 26.800 11.600 27.400 14.600 ;
        RECT 31.600 11.600 32.200 14.600 ;
        RECT 41.200 11.600 41.800 14.600 ;
        RECT 46.000 11.600 46.600 14.600 ;
        RECT 26.800 10.800 28.000 11.600 ;
        RECT 31.600 10.800 32.800 11.600 ;
        RECT 41.200 10.800 42.400 11.600 ;
        RECT 46.000 10.800 47.200 11.600 ;
        RECT 26.800 10.200 27.400 10.800 ;
        RECT 31.600 10.200 32.200 10.800 ;
        RECT 41.200 10.200 41.800 10.800 ;
        RECT 46.000 10.200 46.600 10.800 ;
        RECT 22.200 9.600 24.400 10.200 ;
        RECT 15.600 2.200 16.400 9.600 ;
        RECT 23.600 2.200 24.400 9.600 ;
        RECT 25.200 9.600 27.400 10.200 ;
        RECT 30.000 9.600 32.200 10.200 ;
        RECT 39.600 9.600 41.800 10.200 ;
        RECT 44.400 9.600 46.600 10.200 ;
        RECT 25.200 2.200 26.000 9.600 ;
        RECT 30.000 2.200 30.800 9.600 ;
        RECT 39.600 2.200 40.400 9.600 ;
        RECT 44.400 2.200 45.200 9.600 ;
  END
END dec_to_hex
END LIBRARY

