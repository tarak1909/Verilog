magic
tech scmos
timestamp 1677489954
<< metal1 >>
rect 344 212 392 214
rect 344 208 352 212
rect 356 208 366 212
rect 370 208 380 212
rect 384 208 392 212
rect 344 206 392 208
rect 188 182 196 184
rect 188 178 190 182
rect 194 178 196 182
rect 188 176 196 178
rect 204 182 212 184
rect 204 178 206 182
rect 210 178 212 182
rect 204 176 212 178
rect 284 182 292 184
rect 380 183 388 184
rect 284 178 286 182
rect 290 178 292 182
rect 284 176 292 178
rect 333 182 388 183
rect 333 178 382 182
rect 386 178 388 182
rect 333 177 388 178
rect 380 176 388 177
rect 476 182 484 184
rect 476 178 478 182
rect 482 178 484 182
rect 476 176 484 178
rect 12 162 20 164
rect 12 158 14 162
rect 18 158 20 162
rect 12 156 20 158
rect 60 142 68 144
rect 60 138 62 142
rect 66 138 68 142
rect 60 136 68 138
rect 428 142 436 144
rect 428 138 430 142
rect 434 138 436 142
rect 428 136 436 138
rect 44 122 52 124
rect 44 118 46 122
rect 50 118 52 122
rect 44 116 52 118
rect 92 122 100 124
rect 92 118 94 122
rect 98 118 100 122
rect 92 116 100 118
rect 108 123 116 124
rect 108 122 163 123
rect 108 118 110 122
rect 114 118 163 122
rect 108 117 163 118
rect 236 122 244 124
rect 236 118 238 122
rect 242 118 244 122
rect 108 116 116 117
rect 236 116 244 118
rect 252 122 260 124
rect 252 118 254 122
rect 258 118 260 122
rect 252 116 260 118
rect 300 122 308 124
rect 300 118 302 122
rect 306 118 308 122
rect 300 116 308 118
rect 396 122 404 124
rect 396 118 398 122
rect 402 118 404 122
rect 396 116 404 118
rect 444 122 452 124
rect 444 118 446 122
rect 450 118 452 122
rect 444 116 452 118
rect 104 12 152 14
rect 104 8 112 12
rect 116 8 126 12
rect 130 8 140 12
rect 144 8 152 12
rect 104 6 152 8
<< m2contact >>
rect 352 208 356 212
rect 366 208 370 212
rect 380 208 384 212
rect 190 178 194 182
rect 206 178 210 182
rect 286 178 290 182
rect 382 178 386 182
rect 478 178 482 182
rect 14 158 18 162
rect 62 138 66 142
rect 430 138 434 142
rect 46 118 50 122
rect 94 118 98 122
rect 110 118 114 122
rect 238 118 242 122
rect 254 118 258 122
rect 302 118 306 122
rect 398 118 402 122
rect 446 118 450 122
rect 112 8 116 12
rect 126 8 130 12
rect 140 8 144 12
<< metal2 >>
rect 397 257 435 263
rect 397 243 403 257
rect 28 202 36 204
rect 28 198 30 202
rect 34 198 36 202
rect 28 196 36 198
rect 12 162 20 164
rect 12 158 14 162
rect 18 158 20 162
rect 12 156 20 158
rect 29 163 35 196
rect 45 184 51 243
rect 77 204 83 243
rect 125 204 131 243
rect 76 202 84 204
rect 76 198 78 202
rect 82 198 84 202
rect 76 196 84 198
rect 108 202 116 204
rect 108 198 110 202
rect 114 198 116 202
rect 108 196 116 198
rect 124 202 132 204
rect 124 198 126 202
rect 130 198 132 202
rect 124 196 132 198
rect 44 182 52 184
rect 44 178 46 182
rect 50 178 52 182
rect 44 176 52 178
rect 92 182 100 184
rect 92 178 94 182
rect 98 178 100 182
rect 92 176 100 178
rect 29 157 51 163
rect 45 124 51 157
rect 60 142 68 144
rect 60 138 62 142
rect 66 138 68 142
rect 60 136 68 138
rect 61 124 67 136
rect 93 124 99 176
rect 109 124 115 196
rect 157 184 163 243
rect 237 237 259 243
rect 188 202 196 204
rect 188 198 190 202
rect 194 198 196 202
rect 188 196 196 198
rect 189 184 195 196
rect 156 182 164 184
rect 156 178 158 182
rect 162 178 164 182
rect 156 176 164 178
rect 188 182 196 184
rect 188 178 190 182
rect 194 178 196 182
rect 188 176 196 178
rect 204 182 212 184
rect 204 178 206 182
rect 210 178 212 182
rect 204 176 212 178
rect 237 124 243 237
rect 285 204 291 243
rect 317 237 339 243
rect 365 237 403 243
rect 252 202 260 204
rect 252 198 254 202
rect 258 198 260 202
rect 252 196 260 198
rect 284 202 292 204
rect 284 198 286 202
rect 290 198 292 202
rect 284 196 292 198
rect 253 124 259 196
rect 317 184 323 237
rect 344 212 392 214
rect 344 208 352 212
rect 356 208 366 212
rect 370 208 380 212
rect 384 208 392 212
rect 344 206 392 208
rect 284 182 292 184
rect 284 178 286 182
rect 290 178 292 182
rect 284 176 292 178
rect 316 182 324 184
rect 316 178 318 182
rect 322 178 324 182
rect 316 176 324 178
rect 380 182 388 184
rect 380 178 382 182
rect 386 178 388 182
rect 380 176 388 178
rect 300 162 308 164
rect 300 158 302 162
rect 306 158 308 162
rect 300 156 308 158
rect 301 124 307 156
rect 413 144 419 243
rect 429 204 435 257
rect 477 237 499 243
rect 428 202 436 204
rect 428 198 430 202
rect 434 198 436 202
rect 428 196 436 198
rect 460 202 468 204
rect 460 198 462 202
rect 466 198 468 202
rect 460 196 468 198
rect 461 164 467 196
rect 477 184 483 237
rect 476 182 484 184
rect 476 178 478 182
rect 482 178 484 182
rect 476 176 484 178
rect 460 162 468 164
rect 460 158 462 162
rect 466 158 468 162
rect 460 156 468 158
rect 412 142 420 144
rect 412 138 414 142
rect 418 138 420 142
rect 412 136 420 138
rect 428 142 436 144
rect 428 138 430 142
rect 434 138 436 142
rect 428 136 436 138
rect 444 142 452 144
rect 444 138 446 142
rect 450 138 452 142
rect 444 136 452 138
rect 429 124 435 136
rect 445 124 451 136
rect 44 122 52 124
rect 44 118 46 122
rect 50 118 52 122
rect 44 116 52 118
rect 60 122 68 124
rect 60 118 62 122
rect 66 118 68 122
rect 60 116 68 118
rect 92 122 100 124
rect 92 118 94 122
rect 98 118 100 122
rect 92 116 100 118
rect 108 122 116 124
rect 108 118 110 122
rect 114 118 116 122
rect 108 116 116 118
rect 236 122 244 124
rect 236 118 238 122
rect 242 118 244 122
rect 236 116 244 118
rect 252 122 260 124
rect 252 118 254 122
rect 258 118 260 122
rect 252 116 260 118
rect 300 122 308 124
rect 300 118 302 122
rect 306 118 308 122
rect 300 116 308 118
rect 396 122 404 124
rect 396 118 398 122
rect 402 118 404 122
rect 396 116 404 118
rect 428 122 436 124
rect 428 118 430 122
rect 434 118 436 122
rect 428 116 436 118
rect 444 122 452 124
rect 444 118 446 122
rect 450 118 452 122
rect 444 116 452 118
rect 397 104 403 116
rect 396 102 404 104
rect 396 98 398 102
rect 402 98 404 102
rect 396 96 404 98
rect 104 12 152 14
rect 104 8 112 12
rect 116 8 126 12
rect 130 8 140 12
rect 144 8 152 12
rect 104 6 152 8
<< m3contact >>
rect 30 198 34 202
rect 14 158 18 162
rect 78 198 82 202
rect 110 198 114 202
rect 126 198 130 202
rect 46 178 50 182
rect 94 178 98 182
rect 190 198 194 202
rect 158 178 162 182
rect 206 178 210 182
rect 254 198 258 202
rect 286 198 290 202
rect 352 208 356 212
rect 366 208 370 212
rect 380 208 384 212
rect 286 178 290 182
rect 318 178 322 182
rect 382 178 386 182
rect 302 158 306 162
rect 430 198 434 202
rect 462 198 466 202
rect 462 158 466 162
rect 414 138 418 142
rect 446 138 450 142
rect 62 118 66 122
rect 430 118 434 122
rect 398 98 402 102
rect 112 8 116 12
rect 126 8 130 12
rect 140 8 144 12
<< metal3 >>
rect 344 212 392 216
rect 344 208 350 212
rect 356 208 366 212
rect 370 208 380 212
rect 386 208 392 212
rect 344 204 392 208
rect 28 203 36 204
rect -19 202 36 203
rect -19 198 30 202
rect 34 198 36 202
rect -19 197 36 198
rect 28 196 36 197
rect 76 203 84 204
rect 108 203 116 204
rect 76 202 116 203
rect 76 198 78 202
rect 82 198 110 202
rect 114 198 116 202
rect 76 197 116 198
rect 76 196 84 197
rect 108 196 116 197
rect 124 203 132 204
rect 188 203 196 204
rect 124 202 196 203
rect 124 198 126 202
rect 130 198 190 202
rect 194 198 196 202
rect 124 197 196 198
rect 124 196 132 197
rect 188 196 196 197
rect 252 203 260 204
rect 284 203 292 204
rect 252 202 292 203
rect 252 198 254 202
rect 258 198 286 202
rect 290 198 292 202
rect 252 197 292 198
rect 252 196 260 197
rect 284 196 292 197
rect 428 202 436 204
rect 428 198 430 202
rect 434 198 436 202
rect 428 196 436 198
rect 460 203 468 204
rect 460 202 515 203
rect 460 198 462 202
rect 466 198 515 202
rect 460 197 515 198
rect 460 196 468 197
rect 44 183 52 184
rect 92 183 100 184
rect 44 182 100 183
rect 44 178 46 182
rect 50 178 94 182
rect 98 178 100 182
rect 44 177 100 178
rect 44 176 52 177
rect 92 176 100 177
rect 156 183 164 184
rect 204 183 212 184
rect 156 182 212 183
rect 156 178 158 182
rect 162 178 206 182
rect 210 178 212 182
rect 156 177 212 178
rect 156 176 164 177
rect 204 176 212 177
rect 284 183 292 184
rect 316 183 324 184
rect 284 182 324 183
rect 284 178 286 182
rect 290 178 318 182
rect 322 178 324 182
rect 284 177 324 178
rect 284 176 292 177
rect 316 176 324 177
rect 380 183 388 184
rect 380 182 515 183
rect 380 178 382 182
rect 386 178 515 182
rect 380 177 515 178
rect 380 176 388 177
rect 12 163 20 164
rect -19 162 20 163
rect -19 158 14 162
rect 18 158 20 162
rect -19 157 20 158
rect 12 156 20 157
rect 300 163 308 164
rect 460 163 468 164
rect 300 162 468 163
rect 300 158 302 162
rect 306 158 462 162
rect 466 158 468 162
rect 300 157 468 158
rect 509 157 515 177
rect 300 156 308 157
rect 460 156 468 157
rect 412 143 420 144
rect 444 143 452 144
rect 412 142 452 143
rect 412 138 414 142
rect 418 138 446 142
rect 450 138 452 142
rect 412 137 452 138
rect 412 136 420 137
rect 444 136 452 137
rect 60 123 68 124
rect -19 122 68 123
rect -19 118 62 122
rect 66 118 68 122
rect -19 117 68 118
rect 60 116 68 117
rect 428 123 436 124
rect 428 122 515 123
rect 428 118 430 122
rect 434 118 515 122
rect 428 117 515 118
rect 428 116 436 117
rect 396 103 404 104
rect 428 103 436 104
rect 396 102 436 103
rect 396 98 398 102
rect 402 98 430 102
rect 434 98 436 102
rect 396 97 436 98
rect 396 96 404 97
rect 428 96 436 97
rect 104 12 152 16
rect 104 8 110 12
rect 116 8 126 12
rect 130 8 140 12
rect 146 8 152 12
rect 104 4 152 8
<< m4contact >>
rect 350 208 352 212
rect 352 208 354 212
rect 366 208 370 212
rect 382 208 384 212
rect 384 208 386 212
rect 430 198 434 202
rect 430 98 434 102
rect 110 8 112 12
rect 112 8 114 12
rect 126 8 130 12
rect 142 8 144 12
rect 144 8 146 12
<< metal4 >>
rect 104 12 152 240
rect 104 8 110 12
rect 114 8 126 12
rect 130 8 142 12
rect 146 8 152 12
rect 104 0 152 8
rect 344 212 392 240
rect 344 208 350 212
rect 354 208 366 212
rect 370 208 382 212
rect 386 208 392 212
rect 344 0 392 208
rect 426 202 438 206
rect 426 198 430 202
rect 434 198 438 202
rect 426 102 438 198
rect 426 98 430 102
rect 434 98 438 102
rect 426 94 438 98
use BUFX2  BUFX2_5
timestamp 1677489954
transform -1 0 56 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_7
timestamp 1677489954
transform -1 0 104 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_0_0
timestamp 1677489954
transform 1 0 104 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1677489954
transform 1 0 120 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1677489954
transform 1 0 136 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_1
timestamp 1677489954
transform 1 0 152 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_3
timestamp 1677489954
transform -1 0 248 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_6
timestamp 1677489954
transform 1 0 248 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_8
timestamp 1677489954
transform 1 0 296 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_1_0
timestamp 1677489954
transform 1 0 344 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1677489954
transform 1 0 360 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_2
timestamp 1677489954
transform 1 0 376 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_2
timestamp 1677489954
transform 1 0 392 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_4
timestamp 1677489954
transform 1 0 440 0 -1 210
box -4 -6 52 206
<< labels >>
flabel metal4 s 104 0 152 24 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 344 0 392 24 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 80 240 80 240 7 FreeSans 24 90 0 0 decimal[0]
port 2 nsew
flabel metal2 s 368 240 368 240 3 FreeSans 24 90 0 0 decimal[1]
port 3 nsew
flabel metal2 s 256 240 256 240 3 FreeSans 24 90 0 0 decimal[2]
port 4 nsew
flabel metal2 s 416 240 416 240 3 FreeSans 24 90 0 0 decimal[3]
port 5 nsew
flabel metal3 s -16 200 -16 200 7 FreeSans 24 90 0 0 decimal[4]
port 6 nsew
flabel metal2 s 288 240 288 240 3 FreeSans 24 90 0 0 decimal[5]
port 7 nsew
flabel metal2 s 48 240 48 240 7 FreeSans 24 90 0 0 decimal[6]
port 8 nsew
flabel metal3 s 512 200 512 200 3 FreeSans 24 90 0 0 decimal[7]
port 9 nsew
flabel metal2 s 128 240 128 240 3 FreeSans 24 90 0 0 binary[0]
port 10 nsew
flabel metal3 s 512 120 512 120 3 FreeSans 24 0 0 0 binary[1]
port 11 nsew
flabel metal2 s 160 240 160 240 3 FreeSans 24 90 0 0 binary[2]
port 12 nsew
flabel metal2 s 496 240 496 240 3 FreeSans 24 90 0 0 binary[3]
port 13 nsew
flabel metal3 s -16 160 -16 160 7 FreeSans 24 0 0 0 binary[4]
port 14 nsew
flabel metal2 s 336 240 336 240 3 FreeSans 24 90 0 0 binary[5]
port 15 nsew
flabel metal3 s -16 120 -16 120 7 FreeSans 24 0 0 0 binary[6]
port 16 nsew
flabel metal3 s 512 160 512 160 3 FreeSans 24 0 0 0 binary[7]
port 17 nsew
<< end >>
