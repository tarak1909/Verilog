* NGSPICE file created from dec_to_hex.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

.subckt dec_to_hex vdd gnd decimal[0] decimal[1] decimal[2] decimal[3] decimal[4]
+ decimal[5] decimal[6] decimal[7] hex[0] hex[1] hex[2] hex[3] hex[4] hex[5] hex[6]
+ hex[7]
XFILL_0_0_0 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XFILL_0_0_2 gnd vdd FILL
XBUFX2_1 decimal[0] gnd hex[0] vdd BUFX2
XBUFX2_2 decimal[1] gnd hex[1] vdd BUFX2
XBUFX2_3 decimal[2] gnd hex[2] vdd BUFX2
XBUFX2_4 decimal[3] gnd hex[3] vdd BUFX2
XBUFX2_5 decimal[4] gnd hex[4] vdd BUFX2
XFILL_0_1_0 gnd vdd FILL
XBUFX2_6 decimal[5] gnd hex[5] vdd BUFX2
XFILL_0_1_1 gnd vdd FILL
XBUFX2_7 decimal[6] gnd hex[6] vdd BUFX2
XFILL_0_1_2 gnd vdd FILL
XBUFX2_8 decimal[7] gnd hex[7] vdd BUFX2
.ends

