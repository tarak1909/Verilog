magic
tech scmos
magscale 1 2
timestamp 1677493391
<< metal1 >>
rect 344 206 350 214
rect 358 206 364 214
rect 372 206 378 214
rect 386 206 392 214
rect 333 177 380 183
rect 116 117 163 123
rect 104 6 110 14
rect 118 6 124 14
rect 132 6 138 14
rect 146 6 152 14
<< m2contact >>
rect 350 206 358 214
rect 364 206 372 214
rect 378 206 386 214
rect 188 176 196 184
rect 204 176 212 184
rect 284 176 292 184
rect 380 176 388 184
rect 476 176 484 184
rect 12 156 20 164
rect 60 136 68 144
rect 428 136 436 144
rect 44 116 52 124
rect 92 116 100 124
rect 108 116 116 124
rect 236 116 244 124
rect 252 116 260 124
rect 300 116 308 124
rect 396 116 404 124
rect 444 116 452 124
rect 110 6 118 14
rect 124 6 132 14
rect 138 6 146 14
<< metal2 >>
rect 397 257 435 263
rect 397 243 403 257
rect 29 163 35 196
rect 45 184 51 243
rect 77 204 83 243
rect 125 204 131 243
rect 29 157 51 163
rect 45 124 51 157
rect 61 124 67 136
rect 93 124 99 176
rect 109 124 115 196
rect 157 184 163 243
rect 237 237 259 243
rect 189 184 195 196
rect 237 124 243 237
rect 285 204 291 243
rect 317 237 339 243
rect 365 237 403 243
rect 253 124 259 196
rect 317 184 323 237
rect 344 206 350 214
rect 358 206 364 214
rect 372 206 378 214
rect 386 206 392 214
rect 301 124 307 156
rect 413 144 419 243
rect 429 204 435 257
rect 477 237 499 243
rect 461 164 467 196
rect 477 184 483 237
rect 429 124 435 136
rect 445 124 451 136
rect 397 104 403 116
rect 104 6 110 14
rect 118 6 124 14
rect 132 6 138 14
rect 146 6 152 14
<< m3contact >>
rect 28 196 36 204
rect 12 156 20 164
rect 76 196 84 204
rect 108 196 116 204
rect 124 196 132 204
rect 44 176 52 184
rect 92 176 100 184
rect 188 196 196 204
rect 156 176 164 184
rect 204 176 212 184
rect 252 196 260 204
rect 284 196 292 204
rect 350 206 358 214
rect 364 206 372 214
rect 378 206 386 214
rect 284 176 292 184
rect 316 176 324 184
rect 380 176 388 184
rect 300 156 308 164
rect 428 196 436 204
rect 460 196 468 204
rect 460 156 468 164
rect 412 136 420 144
rect 444 136 452 144
rect 60 116 68 124
rect 428 116 436 124
rect 396 96 404 104
rect 110 6 118 14
rect 124 6 132 14
rect 138 6 146 14
<< metal3 >>
rect 344 214 392 216
rect 344 206 348 214
rect 358 206 364 214
rect 372 206 378 214
rect 388 206 392 214
rect 344 204 392 206
rect -19 197 28 203
rect 84 197 108 203
rect 132 197 188 203
rect 260 197 284 203
rect 468 197 515 203
rect 52 177 92 183
rect 164 177 204 183
rect 292 177 316 183
rect 388 177 515 183
rect -19 157 12 163
rect 308 157 460 163
rect 509 157 515 177
rect 420 137 444 143
rect -19 117 60 123
rect 436 117 515 123
rect 404 97 428 103
rect 104 14 152 16
rect 104 6 108 14
rect 118 6 124 14
rect 132 6 138 14
rect 148 6 152 14
rect 104 4 152 6
<< m4contact >>
rect 348 206 350 214
rect 350 206 356 214
rect 364 206 372 214
rect 380 206 386 214
rect 386 206 388 214
rect 428 196 436 204
rect 428 96 436 104
rect 108 6 110 14
rect 110 6 116 14
rect 124 6 132 14
rect 140 6 146 14
rect 146 6 148 14
<< metal4 >>
rect 104 14 152 240
rect 104 6 108 14
rect 116 6 124 14
rect 132 6 140 14
rect 148 6 152 14
rect 104 0 152 6
rect 344 214 392 240
rect 344 206 348 214
rect 356 206 364 214
rect 372 206 380 214
rect 388 206 392 214
rect 344 0 392 206
rect 426 204 438 206
rect 426 196 428 204
rect 436 196 438 204
rect 426 104 438 196
rect 426 96 428 104
rect 436 96 438 104
rect 426 94 438 96
use BUFX2  BUFX2_5
timestamp 1677493391
transform -1 0 56 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_7
timestamp 1677493391
transform -1 0 104 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_0_0
timestamp 1677493391
transform 1 0 104 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1677493391
transform 1 0 120 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1677493391
transform 1 0 136 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_1
timestamp 1677493391
transform 1 0 152 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_3
timestamp 1677493391
transform -1 0 248 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_6
timestamp 1677493391
transform 1 0 248 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_8
timestamp 1677493391
transform 1 0 296 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_1_0
timestamp 1677493391
transform 1 0 344 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1677493391
transform 1 0 360 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_2
timestamp 1677493391
transform 1 0 376 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_2
timestamp 1677493391
transform 1 0 392 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_4
timestamp 1677493391
transform 1 0 440 0 -1 210
box -4 -6 52 206
<< labels >>
flabel metal4 s 104 0 152 24 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 344 0 392 24 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 80 240 80 240 3 FreeSans 24 90 0 0 decimal[0]
port 2 nsew
flabel metal2 s 368 240 368 240 3 FreeSans 24 90 0 0 decimal[1]
port 3 nsew
flabel metal2 s 256 240 256 240 3 FreeSans 24 90 0 0 decimal[2]
port 4 nsew
flabel metal2 s 416 240 416 240 3 FreeSans 24 90 0 0 decimal[3]
port 5 nsew
flabel metal3 s -16 200 -16 200 7 FreeSans 24 0 0 0 decimal[4]
port 6 nsew
flabel metal2 s 288 240 288 240 3 FreeSans 24 90 0 0 decimal[5]
port 7 nsew
flabel metal2 s 48 240 48 240 3 FreeSans 24 90 0 0 decimal[6]
port 8 nsew
flabel metal3 s 512 200 512 200 3 FreeSans 24 0 0 0 decimal[7]
port 9 nsew
flabel metal2 s 128 240 128 240 3 FreeSans 24 90 0 0 octal[0]
port 10 nsew
flabel metal3 s 512 120 512 120 3 FreeSans 24 0 0 0 octal[1]
port 11 nsew
flabel metal2 s 160 240 160 240 3 FreeSans 24 90 0 0 octal[2]
port 12 nsew
flabel metal2 s 496 240 496 240 3 FreeSans 24 90 0 0 octal[3]
port 13 nsew
flabel metal3 s -16 160 -16 160 7 FreeSans 24 0 0 0 octal[4]
port 14 nsew
flabel metal2 s 336 240 336 240 3 FreeSans 24 90 0 0 octal[5]
port 15 nsew
flabel metal3 s -16 120 -16 120 7 FreeSans 24 0 0 0 octal[6]
port 16 nsew
flabel metal3 s 512 160 512 160 3 FreeSans 24 0 0 0 octal[7]
port 17 nsew
<< end >>
